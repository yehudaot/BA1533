
//`define DEBUG   // in DEBUG mode, we output one bit per clock cycle (useful for faster simulations)

`timescale 1ns/1ns

module async_transmitter(clk, reset_n, TxD_start, TxD_data, TxD, TxD_busy, BaudTick);
input clk, TxD_start, reset_n, BaudTick;
input [7:0] TxD_data;
output TxD, TxD_busy;

parameter RegisterInputData = 1;	// in RegisterInputData mode, the input doesn't have to stay valid while the character is been transmitted

/*
parameter ClkFrequency = 26000000;	// 25MHz
parameter Baud = 115200;

// Baud generator
parameter BaudGeneratorAccWidth = 16;
reg [BaudGeneratorAccWidth:0] BaudGeneratorAcc;
`ifdef DEBUG
wire [BaudGeneratorAccWidth:0] BaudGeneratorInc = 17'h1000;
`else
wire [BaudGeneratorAccWidth:0] BaudGeneratorInc = ((Baud<<(BaudGeneratorAccWidth-4))+(ClkFrequency>>5))/(ClkFrequency>>4);
`endif

wire BaudTick = BaudGeneratorAcc[BaudGeneratorAccWidth];
*/

wire TxD_busy;
//always @(posedge clk) if(TxD_busy) BaudGeneratorAcc <= BaudGeneratorAcc[BaudGeneratorAccWidth-1:0] + BaudGeneratorInc;

// Transmitter state machine
reg [3:0] state;
reg TxD_ready;
//wire TxD_ready = (state==0);
assign TxD_busy = ~TxD_ready;
reg [7:0] TxD_dataReg;
wire [7:0] TxD_dataD = RegisterInputData ? TxD_dataReg : TxD_data;

always @(posedge clk) 
if(TxD_start) 
	TxD_ready <= 1'b0;
else if(BaudTick & (state == 0))
	TxD_ready <= 1'b1;

always @(posedge clk) if(TxD_ready & TxD_start) TxD_dataReg <= TxD_data;
/*
always @ (posedge clk or negedge reset_n)
begin
	if(!reset_n) 
		state <= 4'b0000;
	else if(BaudTick)
	case(state)
		4'b0000: if(TxD_start) state <= 4'b0001;
		4'b0001:  state <= 4'b0100;
		4'b0100:  state <= 4'b1000;  // start
		4'b1000:  state <= 4'b1001;  // bit 0
		4'b1001:  state <= 4'b1010;  // bit 1
		4'b1010:  state <= 4'b1011;  // bit 2
		4'b1011:  state <= 4'b1100;  // bit 3
		4'b1100:  state <= 4'b1101;  // bit 4
		4'b1101:  state <= 4'b1110;  // bit 5
		4'b1110:  state <= 4'b1111;  // bit 6
		4'b1111:  state <= 4'b0010;  // bit 7
		4'b0010:  state <= 4'b0011;  // stop1
		4'b0011:  state <= 4'b0000;  // stop2
		default:  state <= 4'b0000;
	endcase
end
*/

always @ (posedge clk or negedge reset_n)
begin
	if(!reset_n) 
		state <= 4'b0000;
	else if(BaudTick)
	case(state)
		4'b0000: if(TxD_start) state <= 4'b0100;//4'b0001;
		//4'b0001:  state <= 4'b0100;
		4'b0100:  state <= 4'b1000;  // start
		4'b1000:  state <= 4'b1001;  // bit 0
		4'b1001:  state <= 4'b1010;  // bit 1
		4'b1010:  state <= 4'b1011;  // bit 2
		4'b1011:  state <= 4'b1100;  // bit 3
		4'b1100:  state <= 4'b1101;  // bit 4
		4'b1101:  state <= 4'b1110;  // bit 5
		4'b1110:  state <= 4'b1111;  // bit 6
		4'b1111:  state <= 4'b0010;  // bit 7
		4'b0010:  state <= 4'b0000;  // stop1
		//4'b0011:  state <= 4'b0000;  // stop2
		default:  state <= 4'b0000;
	endcase
end

// Output mux
reg muxbit;
always @( * )
case(state[2:0])
	3'd0: muxbit <= TxD_dataD[0];
	3'd1: muxbit <= TxD_dataD[1];
	3'd2: muxbit <= TxD_dataD[2];
	3'd3: muxbit <= TxD_dataD[3];
	3'd4: muxbit <= TxD_dataD[4];
	3'd5: muxbit <= TxD_dataD[5];
	3'd6: muxbit <= TxD_dataD[6];
	3'd7: muxbit <= TxD_dataD[7];
endcase

// Put together the start, data and stop bits
reg TxD;
always @(posedge clk) TxD <= (state<4) | (state[3] & muxbit);  // register the output to make it glitch free

endmodule
